/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� DDS.v
** �������ڣ�
** ����������DDS�źŷ�����Ƕ��ʽ�߼������ǵĵ���
** Ӳ��ƽ̨�������ϵ�һ��������
** ��Ȩ������������������֪ʶ��Ȩ,�������������ѧϰ.
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module DDS(
			clk,
			dds_data_out,
			set_waveform,
			set_f,
			set_a,
			set_p
          );
input         clk;//ʱ������
input  [1:0]  set_waveform;
input  [20:0] set_f;
input  [4:0]  set_a;
input  [8:0]  set_p;
output [9:0]  dds_data_out;

wire          clk;
wire   [1:0]  set_waveform;
wire   [20:0] set_f;
wire   [4:0]  set_a;
wire   [9:0]  set_p;
wire   [9:0]  dds_data_out;
/**************������***************/
wire   [31:0] f32_bus;//ACƵ�ʿ���������
wire   [31:0] reg32_out;//32λ�Ĵ������
wire   [31:0] reg32_in;//32λ�Ĵ�������
wire   [8:0]  reg10_in;
wire   [8:0]  reg10_out_address;
/**************����Ĵ���******************/
wire   [9:0]  sin_data;
wire   [9:0]  tri_data;
wire   [9:0]  squ_data;
//wire   [9:0]  saw_data;
reg    [9:0]  dds_data_reg; 
reg    [20:0] set_f_reg;     
/***********************************/
assign f32_bus[31:21]=11'b000_0000_0000;//��ʼ��,��λ�õ�
assign f32_bus[20:0]=set_f_reg;    //��λ��������DDS�����Ƶ��
/*********************Ԫ������************************************/
       adder_32 u1(.data1(f32_bus),.data2(reg32_out),.sum(reg32_in));
       reg32    u2(.clk(clk),.data_in(reg32_in),.data_out(reg32_out));
       adder_10 u7(.data1(set_p),.data2(reg32_out[31:23]),.sum(reg10_in));
       reg_10   u8(.clk(clk),.data_in(reg10_in),.data_out(reg10_out_address));
/*****************����ѡ��*******************************************/
       sin_rom  u3(.address(reg10_out_address),.clock(clk),.q(sin_data));//����
       tri_rom  u4(.address(reg10_out_address),.clock(clk),.q(tri_data));
       squ_rom  u5(.address(reg10_out_address),.clock(clk),.q(squ_data));
//       saw_rom  u6(.address(reg10_out_address),.clock(clk),.q(saw_data));
/***********************���ò��κ�����Ƶ��***************************/
    always @(set_waveform,sin_data,tri_data,squ_data)
      begin 
        case (set_waveform)
          2'b00://���Ҳ�
               begin 
                 dds_data_reg<=sin_data; 
                 set_f_reg<=set_f;//���÷�ΧΪ100Hz��20KHz
               end
          2'b01://���ǲ�
               begin
                 dds_data_reg<=tri_data;
                 set_f_reg<=21'd85899;//�̶�Ϊ1KHz
               end
          2'b10:
               begin
                 dds_data_reg<=squ_data;//����
                 set_f_reg<=21'd85899;//�̶�Ϊ1KHz
               end
        default:
               begin
                  dds_data_reg<=sin_data;//���Ҳ�
                  set_f_reg<=set_f;//���÷�ΧΪ100Hz��20KHz
               end
        endcase;
      end 
/***********************���õ�ѹ��ֵ***************************/
assign dds_data_out=dds_data_reg*3/10;//���õ�ѹ��ֵ
endmodule





