/********************************��Ȩ����**************************************
**                              �������Ŷ�
**                            
**----------------------------�ļ���Ϣ--------------------------
** �ļ����ƣ� adder_10.v
** ����������10λ�ۼ���
**---------------------------�޸��ļ��������Ϣ----------------
** �޸��ˣ�
** �޸����ڣ�		
** �޸����ݣ�
*******************************************************************************/
module adder_10(
                data1,
                data2,
                sum);
input [8:0] data1,data2;//������1��2
output [8:0] sum;//�����

wire [8:0] data1,data2;
wire [8:0] sum;

assign sum=data1+data2;

endmodule
